LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

PACKAGE array32 IS
    TYPE array32bits32 IS ARRAY (0 TO 31) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
END PACKAGE array32;